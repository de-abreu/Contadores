-- Copyright (C) 2021  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- PROGRAM		"Quartus Prime"
-- VERSION		"Version 21.1.0 Build 842 10/21/2021 SJ Lite Edition"
-- CREATED		"Tue Sep 17 17:36:30 2024"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY Rotate IS 
	PORT
	(
		Clock :  IN  STD_LOGIC;
		set :  IN  STD_LOGIC;
		h00 :  OUT  STD_LOGIC;
		h01 :  OUT  STD_LOGIC;
		h02 :  OUT  STD_LOGIC;
		h03 :  OUT  STD_LOGIC;
		h04 :  OUT  STD_LOGIC;
		h05 :  OUT  STD_LOGIC;
		h06 :  OUT  STD_LOGIC;
		h10 :  OUT  STD_LOGIC;
		h11 :  OUT  STD_LOGIC;
		h12 :  OUT  STD_LOGIC;
		h13 :  OUT  STD_LOGIC;
		h14 :  OUT  STD_LOGIC;
		h15 :  OUT  STD_LOGIC;
		h16 :  OUT  STD_LOGIC;
		h20 :  OUT  STD_LOGIC;
		h21 :  OUT  STD_LOGIC;
		h22 :  OUT  STD_LOGIC;
		h23 :  OUT  STD_LOGIC;
		h24 :  OUT  STD_LOGIC;
		h25 :  OUT  STD_LOGIC;
		h26 :  OUT  STD_LOGIC
	);
END Rotate;

ARCHITECTURE bdf_type OF Rotate IS 

COMPONENT \4bit_d_flipflop\
	PORT(p3 : IN STD_LOGIC;
		 p2 : IN STD_LOGIC;
		 p1 : IN STD_LOGIC;
		 p0 : IN STD_LOGIC;
		 Clk : IN STD_LOGIC;
		 Clear : IN STD_LOGIC;
		 n3 : OUT STD_LOGIC;
		 n2 : OUT STD_LOGIC;
		 n1 : OUT STD_LOGIC;
		 n0 : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT hexdisplay
	PORT(x3 : IN STD_LOGIC;
		 x2 : IN STD_LOGIC;
		 x1 : IN STD_LOGIC;
		 x0 : IN STD_LOGIC;
		 h0 : OUT STD_LOGIC;
		 h1 : OUT STD_LOGIC;
		 h2 : OUT STD_LOGIC;
		 h3 : OUT STD_LOGIC;
		 h4 : OUT STD_LOGIC;
		 h5 : OUT STD_LOGIC;
		 h6 : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT \4bit_multiplexer\
	PORT(i31 : IN STD_LOGIC;
		 i30 : IN STD_LOGIC;
		 i21 : IN STD_LOGIC;
		 i20 : IN STD_LOGIC;
		 i11 : IN STD_LOGIC;
		 i10 : IN STD_LOGIC;
		 i01 : IN STD_LOGIC;
		 i00 : IN STD_LOGIC;
		 selection : IN STD_LOGIC;
		 o3 : OUT STD_LOGIC;
		 o2 : OUT STD_LOGIC;
		 o1 : OUT STD_LOGIC;
		 o0 : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT \2\
	PORT(		 d3 : OUT STD_LOGIC;
		 d2 : OUT STD_LOGIC;
		 d1 : OUT STD_LOGIC;
		 d0 : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT e
	PORT(		 d3 : OUT STD_LOGIC;
		 d2 : OUT STD_LOGIC;
		 d1 : OUT STD_LOGIC;
		 d0 : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT d
	PORT(		 d3 : OUT STD_LOGIC;
		 d2 : OUT STD_LOGIC;
		 d1 : OUT STD_LOGIC;
		 d0 : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT rotation
	PORT(p3 : IN STD_LOGIC;
		 p2 : IN STD_LOGIC;
		 p1 : IN STD_LOGIC;
		 p0 : IN STD_LOGIC;
		 n3 : OUT STD_LOGIC;
		 n2 : OUT STD_LOGIC;
		 n1 : OUT STD_LOGIC;
		 n0 : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	clk :  STD_LOGIC;
SIGNAL	s :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_60 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_61 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_62 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_63 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_64 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_65 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_66 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_67 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_68 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_69 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_70 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_71 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_35 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_37 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_39 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_43 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_45 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_47 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_48 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_49 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_50 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_51 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_52 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_53 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_54 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_55 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_56 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_57 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_58 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_59 :  STD_LOGIC;


BEGIN 



b2v_ff0 : \4bit_d_flipflop\
PORT MAP(p3 => SYNTHESIZED_WIRE_0,
		 p2 => SYNTHESIZED_WIRE_1,
		 p1 => SYNTHESIZED_WIRE_2,
		 p0 => SYNTHESIZED_WIRE_3,
		 Clk => clk,
		 n3 => SYNTHESIZED_WIRE_48,
		 n2 => SYNTHESIZED_WIRE_49,
		 n1 => SYNTHESIZED_WIRE_50,
		 n0 => SYNTHESIZED_WIRE_51);


b2v_ff1 : \4bit_d_flipflop\
PORT MAP(p3 => SYNTHESIZED_WIRE_4,
		 p2 => SYNTHESIZED_WIRE_5,
		 p1 => SYNTHESIZED_WIRE_6,
		 p0 => SYNTHESIZED_WIRE_7,
		 Clk => clk,
		 n3 => SYNTHESIZED_WIRE_52,
		 n2 => SYNTHESIZED_WIRE_53,
		 n1 => SYNTHESIZED_WIRE_54,
		 n0 => SYNTHESIZED_WIRE_55);


b2v_ff2 : \4bit_d_flipflop\
PORT MAP(p3 => SYNTHESIZED_WIRE_8,
		 p2 => SYNTHESIZED_WIRE_9,
		 p1 => SYNTHESIZED_WIRE_10,
		 p0 => SYNTHESIZED_WIRE_11,
		 Clk => clk,
		 n3 => SYNTHESIZED_WIRE_56,
		 n2 => SYNTHESIZED_WIRE_57,
		 n1 => SYNTHESIZED_WIRE_58,
		 n0 => SYNTHESIZED_WIRE_59);


b2v_hex0 : hexdisplay
PORT MAP(x3 => SYNTHESIZED_WIRE_60,
		 x2 => SYNTHESIZED_WIRE_61,
		 x1 => SYNTHESIZED_WIRE_62,
		 x0 => SYNTHESIZED_WIRE_63,
		 h0 => h00,
		 h1 => h01,
		 h2 => h02,
		 h3 => h03,
		 h4 => h04,
		 h5 => h05,
		 h6 => h06);


b2v_hex1 : hexdisplay
PORT MAP(x3 => SYNTHESIZED_WIRE_64,
		 x2 => SYNTHESIZED_WIRE_65,
		 x1 => SYNTHESIZED_WIRE_66,
		 x0 => SYNTHESIZED_WIRE_67,
		 h0 => h10,
		 h1 => h11,
		 h2 => h12,
		 h3 => h13,
		 h4 => h14,
		 h5 => h15,
		 h6 => h16);


b2v_hex2 : hexdisplay
PORT MAP(x3 => SYNTHESIZED_WIRE_68,
		 x2 => SYNTHESIZED_WIRE_69,
		 x1 => SYNTHESIZED_WIRE_70,
		 x0 => SYNTHESIZED_WIRE_71,
		 h0 => h20,
		 h1 => h21,
		 h2 => h22,
		 h3 => h23,
		 h4 => h24,
		 h5 => h25,
		 h6 => h26);


b2v_inst : \4bit_multiplexer\
PORT MAP(i31 => SYNTHESIZED_WIRE_68,
		 i30 => SYNTHESIZED_WIRE_25,
		 i21 => SYNTHESIZED_WIRE_69,
		 i20 => SYNTHESIZED_WIRE_27,
		 i11 => SYNTHESIZED_WIRE_70,
		 i10 => SYNTHESIZED_WIRE_29,
		 i01 => SYNTHESIZED_WIRE_71,
		 i00 => SYNTHESIZED_WIRE_31,
		 selection => s,
		 o3 => SYNTHESIZED_WIRE_8,
		 o2 => SYNTHESIZED_WIRE_9,
		 o1 => SYNTHESIZED_WIRE_10,
		 o0 => SYNTHESIZED_WIRE_11);


b2v_inst1 : \4bit_multiplexer\
PORT MAP(i31 => SYNTHESIZED_WIRE_64,
		 i30 => SYNTHESIZED_WIRE_33,
		 i21 => SYNTHESIZED_WIRE_65,
		 i20 => SYNTHESIZED_WIRE_35,
		 i11 => SYNTHESIZED_WIRE_66,
		 i10 => SYNTHESIZED_WIRE_37,
		 i01 => SYNTHESIZED_WIRE_67,
		 i00 => SYNTHESIZED_WIRE_39,
		 selection => s,
		 o3 => SYNTHESIZED_WIRE_4,
		 o2 => SYNTHESIZED_WIRE_5,
		 o1 => SYNTHESIZED_WIRE_6,
		 o0 => SYNTHESIZED_WIRE_7);


b2v_inst2 : \4bit_multiplexer\
PORT MAP(i31 => SYNTHESIZED_WIRE_60,
		 i30 => SYNTHESIZED_WIRE_41,
		 i21 => SYNTHESIZED_WIRE_61,
		 i20 => SYNTHESIZED_WIRE_43,
		 i11 => SYNTHESIZED_WIRE_62,
		 i10 => SYNTHESIZED_WIRE_45,
		 i01 => SYNTHESIZED_WIRE_63,
		 i00 => SYNTHESIZED_WIRE_47,
		 selection => s,
		 o3 => SYNTHESIZED_WIRE_0,
		 o2 => SYNTHESIZED_WIRE_1,
		 o1 => SYNTHESIZED_WIRE_2,
		 o0 => SYNTHESIZED_WIRE_3);


b2v_preset0 : \2\
PORT MAP(		 d3 => SYNTHESIZED_WIRE_41,
		 d2 => SYNTHESIZED_WIRE_43,
		 d1 => SYNTHESIZED_WIRE_45,
		 d0 => SYNTHESIZED_WIRE_47);


b2v_preset1 : e
PORT MAP(		 d3 => SYNTHESIZED_WIRE_33,
		 d2 => SYNTHESIZED_WIRE_35,
		 d1 => SYNTHESIZED_WIRE_37,
		 d0 => SYNTHESIZED_WIRE_39);


b2v_preset2 : d
PORT MAP(		 d3 => SYNTHESIZED_WIRE_25,
		 d2 => SYNTHESIZED_WIRE_27,
		 d1 => SYNTHESIZED_WIRE_29,
		 d0 => SYNTHESIZED_WIRE_31);


b2v_rot0 : rotation
PORT MAP(p3 => SYNTHESIZED_WIRE_48,
		 p2 => SYNTHESIZED_WIRE_49,
		 p1 => SYNTHESIZED_WIRE_50,
		 p0 => SYNTHESIZED_WIRE_51,
		 n3 => SYNTHESIZED_WIRE_60,
		 n2 => SYNTHESIZED_WIRE_61,
		 n1 => SYNTHESIZED_WIRE_62,
		 n0 => SYNTHESIZED_WIRE_63);


b2v_rot1 : rotation
PORT MAP(p3 => SYNTHESIZED_WIRE_52,
		 p2 => SYNTHESIZED_WIRE_53,
		 p1 => SYNTHESIZED_WIRE_54,
		 p0 => SYNTHESIZED_WIRE_55,
		 n3 => SYNTHESIZED_WIRE_64,
		 n2 => SYNTHESIZED_WIRE_65,
		 n1 => SYNTHESIZED_WIRE_66,
		 n0 => SYNTHESIZED_WIRE_67);


b2v_rot2 : rotation
PORT MAP(p3 => SYNTHESIZED_WIRE_56,
		 p2 => SYNTHESIZED_WIRE_57,
		 p1 => SYNTHESIZED_WIRE_58,
		 p0 => SYNTHESIZED_WIRE_59,
		 n3 => SYNTHESIZED_WIRE_68,
		 n2 => SYNTHESIZED_WIRE_69,
		 n1 => SYNTHESIZED_WIRE_70,
		 n0 => SYNTHESIZED_WIRE_71);

s <= set;
clk <= Clock;

END bdf_type;